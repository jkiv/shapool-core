`define TARGET 34
