`define TARGET 39
