`define TARGET 33
