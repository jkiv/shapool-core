`define TARGET 35
