`define TARGET 36
