`define TARGET 40
