`define TARGET 32
