`define TARGET 44
