`define TARGET 42
