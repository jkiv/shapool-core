`define TARGET 37
