`define TARGET 43
