`define TARGET 45
