`define TARGET 41
