`define TARGET 38
